module datapath()